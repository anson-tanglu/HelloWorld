class test; 
/**
* @brief new
*
*/
function new()
begin
	printf("ok");	
end
endclass
